program main;
  initial forever $display("SPAM");
endprogram
