-- Single line commment in VHDL
